module check(output a,output c,output d,output e,output f,output g,output h,output j,output k,output l,output m,output p,output r,output s,output t,output u,output w,output x,output y,output z,output q1,output w1,output e1,output r1,output t1,output y1,output u1,output i1,output o1,output p1,output a1,output s1,output d1,output f1,output g1,output h1,output j1,output l2,output k1,output l1);
assign { a,c,d,e,f,g,h,j,k,l,m,p,r,s,t,u,w,x,y,z,q1,w1,e1,r1,t1,y1,u1,i1,o1,p1,a1,s1,d1,f1,g1,h1,j1,k1,l1,l2} = 46'b1111111111111111111111111111111111111111111111;
endmodule
