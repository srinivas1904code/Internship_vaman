// write a simple verilog program that implement 
module hello(y,x);
output y;
input x;
assign y =!x;
endmodule
